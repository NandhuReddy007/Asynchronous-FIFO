package pkg;

  int no_txn=20;
  `include "transactor.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "receiver.sv"
  `include "scoreboard.sv"
  `include "environment.sv"


endpackage
