class transactor;
  
  rand bit[7:0] d_in;

endclass
